// - - - - - UVM TESTBENCH FOR DECODE UNIT OF RISC-V CORE - - - - - //

// - - - - - TRANSACTION - - - - - //
//

