`ifndef OPCODES_SVH
`define OPCODES_SVH

parameter I_TYPE_OPCODE = 7'b0000011;
