// - - - - - IMMEDIATE GENERATOR - - - - - //
module immediate_gen (
    input [6:0] i_opcode,
    input [31:0] i_instr,
    output [31:0] o_ext_imm
);


endmodule